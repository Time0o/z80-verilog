localparam OP_PREFIX_NONE  = 7'h00;
localparam OP_PREFIX_DD    = 7'h03;
localparam OP_PREFIX_FD    = 7'h05;
localparam OP_PREFIX_ED    = 7'h09;
localparam OP_PREFIX_CB    = 7'h11;
localparam OP_PREFIX_DD_CB = 7'h21;
localparam OP_PREFIX_FD_CB = 7'h41;
