`include "alu.vh"
`include "fsm.vh"
`include "interrupt.vh"
`include "opcode.vh"
`include "regfile.vh"
