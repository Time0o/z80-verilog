localparam FLAG_IDX_S  = 5;
localparam FLAG_IDX_Z  = 4;
localparam FLAG_IDX_H  = 3;
localparam FLAG_IDX_PV = 2;
localparam FLAG_IDX_N  = 1;
localparam FLAG_IDX_C  = 0;
