/*****************************************************************************
 Processor State
 *****************************************************************************/
`define OP_PREFIX_WIDTH 7
`define FSM_STATE_WIDTH 46
`define INT_MODE_WIDTH 2

/*****************************************************************************
 Muxing
 *****************************************************************************/
`define MUX_ALU_OP_A_SEL_WIDTH 5
`define MUX_ALU_OP_B_SEL_WIDTH 4
`define MUX_INT_BUS_SEL_WIDTH 7
`define MUX_MEM_ADDR_SEL_WIDTH 6
`define MUX_MEM_DOUT_SEL_WIDTH 6

/*****************************************************************************
 Register File
 *****************************************************************************/
`define REG_SELECT_8BIT_WIDTH 7
`define REG_SELECT_16BIT_WIDTH 7
`define REG_SELECT_WIDTH 14

/*****************************************************************************
 ALU
 *****************************************************************************/
`define ALU_MODE_WIDTH 37
