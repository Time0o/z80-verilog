localparam ALU_MODE_ADD       = 37'h0000000000;
localparam ALU_MODE_ADC       = 37'h0000000001;
localparam ALU_MODE_SUB       = 37'h0000000002;
localparam ALU_MODE_SBC       = 37'h0000000004;
localparam ALU_MODE_ADD_16BIT = 37'h0000000008;
localparam ALU_MODE_ADC_16BIT = 37'h0000000010;
localparam ALU_MODE_SBC_16BIT = 37'h0000000020;
localparam ALU_MODE_AND       = 37'h0000000040;
localparam ALU_MODE_OR        = 37'h0000000080;
localparam ALU_MODE_XOR       = 37'h0000000100;
localparam ALU_MODE_CP        = 37'h0000000200;
localparam ALU_MODE_INC       = 37'h0000000400;
localparam ALU_MODE_DEC       = 37'h0000000800;
localparam ALU_MODE_CPL       = 37'h0000001000;
localparam ALU_MODE_NEG       = 37'h0000002000;
localparam ALU_MODE_CCF       = 37'h0000004000;
localparam ALU_MODE_SCF       = 37'h0000008000;
localparam ALU_MODE_RLCA      = 37'h0000010000;
localparam ALU_MODE_RLA       = 37'h0000020000;
localparam ALU_MODE_RRCA      = 37'h0000040000;
localparam ALU_MODE_RRA       = 37'h0000080000;
localparam ALU_MODE_RLC       = 37'h0000100000;
localparam ALU_MODE_RL        = 37'h0000200000;
localparam ALU_MODE_RRC       = 37'h0000400000;
localparam ALU_MODE_RR        = 37'h0000800000;
localparam ALU_MODE_SLA       = 37'h0001000000;
localparam ALU_MODE_SRA       = 37'h0002000000;
localparam ALU_MODE_SRL       = 37'h0004000000;
localparam ALU_MODE_RLD       = 37'h0008000000;
localparam ALU_MODE_RRD       = 37'h0010000000;
localparam ALU_MODE_BIT       = 37'h0020000000;
localparam ALU_MODE_SET       = 37'h0040000000;
localparam ALU_MODE_RES       = 37'h0080000000;
localparam ALU_MODE_IN        = 37'h0100000000;
localparam ALU_MODE_INI       = 37'h0200000000;
localparam ALU_MODE_LDAI      = 37'h0400000000;
localparam ALU_MODE_CPB       = 37'h0800000000;
localparam ALU_MODE_DAA       = 37'h1000000000;
