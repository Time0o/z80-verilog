localparam INT_MODE_0 = 2'b00;
localparam INT_MODE_1 = 2'b01;
localparam INT_MODE_2 = 2'b10;
